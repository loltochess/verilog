module betting();

endmodule
