module bet_controller(clk,nRST,state,clr,player1_en,player2_en,player1_raise,player1_call,player2_raise,player2_call);


endmodule
